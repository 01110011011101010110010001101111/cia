module video_sig_gen
#(
  parameter ACTIVE_H_PIXELS = 1280,
  parameter H_FRONT_PORCH = 110,
  parameter H_SYNC_WIDTH = 40,
  parameter H_BACK_PORCH = 220,
  parameter ACTIVE_LINES = 720,
  parameter V_FRONT_PORCH = 5,
  parameter V_SYNC_WIDTH = 5,
  parameter V_BACK_PORCH = 20,
  parameter FPS = 60)
(
  input wire pixel_clk_in,
  input wire rst_in,
  output logic [$clog2(TOTAL_PIXELS)-1:0] hcount_out,
  output logic [$clog2(TOTAL_LINES)-1:0] vcount_out,
  output logic vs_out, //vertical sync out
  output logic hs_out, //horizontal sync out
  output logic ad_out,
  output logic nf_out, //single cycle enable signal
  output logic [5:0] fc_out); //frame

  localparam TOTAL_PIXELS = (ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH + H_BACK_PORCH); // * (V_FRONT_PORCH + ACTIVE_LINES + V_SYNC_WIDTH + V_BACK_PORCH); //figure this out
  localparam TOTAL_LINES = (V_FRONT_PORCH + ACTIVE_LINES + V_SYNC_WIDTH + V_BACK_PORCH); //figure this out

  logic rst_down = 0;
  always_ff @(posedge pixel_clk_in) begin
    if (rst_in) begin
        rst_down <= 1;
        ad_out <= 0;
        hs_out <= 0;
        vs_out <= 0;
        fc_out <= 0;
        nf_out <= 0;
        hcount_out <= 0;
        vcount_out <= 0;
    end else if (rst_down) begin
        rst_down <= 0;
        hcount_out <= 0;
        vcount_out <= 0;
        ad_out <= 1;
    end else begin
        // update ad_out (and account for wraparound)
        if (
            // we're at the edges
            (hcount_out+1 < ACTIVE_H_PIXELS || hcount_out + 1 == TOTAL_PIXELS) && 
            (
                // if we're within ACTIVE_LINES (when we're not about to increment vcount_out)
                (vcount_out < ACTIVE_LINES && hcount_out + 1 != TOTAL_PIXELS) || 
                // if we're within or at 0 when we're about to increment vcount_out
                ((vcount_out + 1 < ACTIVE_LINES || vcount_out + 1 == TOTAL_LINES) && hcount_out + 1 == TOTAL_PIXELS)
            )
        ) begin
            ad_out <= 1;
        end else begin
            ad_out <= 0;
        end

        // update hs_out
        if (ACTIVE_H_PIXELS + H_FRONT_PORCH <= hcount_out + 1 && hcount_out + 1 < ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH) begin
            hs_out <= 1;
        end else begin
            hs_out <= 0;
        end 

        // update the counts
        if (hcount_out + 1 == TOTAL_PIXELS) begin
            vcount_out <= vcount_out == TOTAL_LINES - 1 ? 0 : vcount_out + 1; 

            // update vs_out
            if (ACTIVE_LINES + V_FRONT_PORCH <= vcount_out + 1 && vcount_out + 1 < ACTIVE_LINES + V_FRONT_PORCH + V_SYNC_WIDTH) begin
                vs_out <= 1;
            end else begin
                vs_out <= 0;
            end 

        end
        hcount_out <= hcount_out == TOTAL_PIXELS - 1 ? 0 : hcount_out + 1; 

        // update fc_out + nf_out
        // NOTE: may need to offset by 1
        if (vcount_out == ACTIVE_LINES && hcount_out + 1 == ACTIVE_H_PIXELS) begin
            fc_out <= fc_out == FPS-1 ? 0 : fc_out + 1;
            nf_out <= 1;
        end else begin
            nf_out <= 0;
        end



    end
  end


  //your code here


endmodule
